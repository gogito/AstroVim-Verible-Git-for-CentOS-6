package pkg;
  import uvm_pkg::*;
  
  `include "uvm_macros.svh"
  `include "sequence_item.sv"
  `include "sequence.sv"
  `include "other_sequence.sv"
  `include "monitor.sv"
  `include "driver.sv"
  `include "scoreboard.sv"
  `include "agent.sv"
  `include "env.sv"
  `include "test.sv"
endpackage